module info