module apache

