module info

pub struct HW {
	
}