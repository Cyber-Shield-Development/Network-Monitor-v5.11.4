module config 

pub struct ProtectionSettings 
{
	
}