module nginx
