module nginx

