module info

