module shield

pub const (
	ssh_protocol = ""
	openvpn_protocol = ""
	apache_protocol = ""
)

pub fn parse_incoming_request(request_info string, pkt_data string) 
{

}